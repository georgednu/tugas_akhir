//`define WIDTH 32
//`define FRAC 20

`define N_MAX 6
`define RK_ORD 4
//`define RK_ORD_3
//`define RK_ORD_2
//`define RK_ORD_1

`define CLK_COUNTER 25 //2MHz clock counter for 50MHz
//`define time_step 2147 //Approx 200kHz/

`define DMA_WIDTH 64
`define PARAMETER_WIDTH 43
`define PARAMETER_FRAC 32
`define STATE_WIDTH 43
`define STATE_FRAC 32